/*
    //------------------------------------------------------------------------------------
    //      Генератор одиночного импульса заданной длительности после подачи питания
    initialpulse
    #(
        .LEN    (), // Длительность импульса
        .POL    ()  // Активный уровень импульса
    )
    the_initialpulse
    (
        // Тактирование
        .clk    (), // i
        
        // Импульс, генерируемый при старте
        .pulse  ()  // o
    ); // the_initialpulse
*/

module initialpulse
#(
    parameter int unsigned  LEN = 10,   // Длительность импульса (от первого фронта clk)
    parameter logic         POL = 1'b1  // Активный уровень импульса
)
(
    // Тактирование
    input  logic            clk,
    
    // Импульс, генерируемый при старте
    output logic            pulse
);
    //------------------------------------------------------------------------------------
    //      Описание констант
    localparam int unsigned CWIDTH = LEN < 1 ? 1 : $clog2(LEN + 1);
    
    //------------------------------------------------------------------------------------
    //      Объявление сигналов
    logic [CWIDTH - 1 : 0]  delay_cnt;
    logic                   pulse_reg;
    
    //------------------------------------------------------------------------------------
    //      Счетчик задержки
    initial delay_cnt = LEN[CWIDTH - 1 : 0];
    always @(posedge clk)
        delay_cnt <= delay_cnt - (delay_cnt != 0);
    
    //------------------------------------------------------------------------------------
    //      Регистр генерируемого импульса
    initial pulse_reg = POL;
    always @(posedge clk)
        pulse_reg <= (LEN == 0) ? ~POL : (delay_cnt != 0) ^ (~POL);
    assign pulse = pulse_reg;
    
endmodule: initialpulse