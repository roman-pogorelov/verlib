/****************************************************************************************
*                                                                                       *
* clockmon                                                                              *
*                                                                                       *
* Модуль контроля тактового сигнала.                                                    *
*                                                                                       *
*       Модуль выполняет контроль наличия тактового сигнала monclk по опорному          *
* тактовому сигналу refclk. При обнаружении стабильных изменений на входе monclk        *
* признак наличия detected устанавливается, при их пропадании - сбрасывается.           *
*                                                                                       *
*   Параметры модуля:                                                                   *
*       FREQRATIO - отношение частоты опорного сигнала к частоте контролируемого,       *
*       округленное до ближайшего большего, т.е.                                        *
*                   FREQRATIO = ceil(FREQ(refclk)/FREQ(monclk)).                        *
*       В случае, если на вход monclk предполагается подавать сигнал, частота которого  *
*       в процессе работы может меняться в некотором диапазоне, то для расчета          *
*       FREQRATIO необходимо использовать МИНИМАЛЬНОЕ значение диапазона.               *
*                                                                                       *
*****************************************************************************************
* Создан:                                                                               *
*       Погорелов Р.А., подр. 171, 2015.12.29                                           *
*                                                                                       *
* Изменения:                                                                            *
*                                                                                       *
*****************************************************************************************
* Необходимые изменения:                                                                *
*                                                                                       *
****************************************************************************************/

/*
    //------------------------------------------------------------------------------------
    //      Модуль контроля тактового сигнала
    clockmon
    #(
       .FREQRATIO   ()  // FREQRATIO = ceil(FREQ(refclk)/FREQ(monclk))
    )
    the_clockmon
    (
        // Общий асинхронный сброс
        .reset      (), // i
        
        // Контролируемый тактовый сигнал
        .monclk     (), // i
        
        // Опорный (стабильный) тактовый сигнал
        .refclk     (), // i
        
        // Признак наличия контролируемого 
        // тактового сигнала
        .detected   ()  // o
    ); // the_clockmon
*/
module clockmon
#(
    parameter int unsigned  FREQRATIO = 2   // FREQRATIO = ceil(FREQ(monclk)/FREQ(refclk))
)
(
    // Общий асинхронный сброс
    input  logic            reset,
    
    // Контролируемый тактовый сигнал
    input  logic            monclk,
    
    // Опорный (стабильный) тактовый сигнал
    input  logic            refclk,
    
    // Признак наличия контролируемого 
    // тактового сигнала
    output logic            detected
);
    //------------------------------------------------------------------------------------
    //      Длина регистровых ступеней
    localparam CYCLES = 3;
    
    //------------------------------------------------------------------------------------
    //      Количество дополнительных тактов для перестраховки с учетом метастабильности
    localparam ADDCYCLES = 2;
    
    //------------------------------------------------------------------------------------
    //      Количество тактов частоты refclk, в течение которых гарантированно должен
    //      быть сформирован хотябы один импульс
    localparam COUNT = (CYCLES + ADDCYCLES)*(1 + FREQRATIO);
    
    //------------------------------------------------------------------------------------
    //      Разрядность счетчика обнаружения
    localparam CWIDTH = $clog2(COUNT);
    
    //------------------------------------------------------------------------------------
    //      Максимальное значение счетчика обнаружения
    localparam logic [CWIDTH - 1 : 0] CMAX = COUNT[CWIDTH - 1 : 0] - 1'b1;
    
    //------------------------------------------------------------------------------------
    //      Описание сигналов
    logic                   pulse_reg;      // Регистр импульсов наличия контролируемого тактового сигнала
    logic [CWIDTH - 1 : 0]  detect_cnt;     // Счетчик обнаружения
    logic                   detect_reg;     // Регистр обнаружения
    
    //------------------------------------------------------------------------------------
    //      Объявление сигналов с учетом требований синтеза и проверки Altera
    (*altera_attribute = "-name SDC_STATEMENT \"set_false_path -from [get_registers {*clockmon:*|mon_reg[*]}] -to [get_registers {*clockmon:*|ref_reg[*]}]\""*) reg [CYCLES - 1 : 0] ref_reg;
    (*altera_attribute = "-name SDC_STATEMENT \"set_false_path -from [get_registers {*clockmon:*|ref_reg[*]}] -to [get_registers {*clockmon:*|mon_reg[*]}]\""*) reg [CYCLES - 1 : 0] mon_reg;
    
    //------------------------------------------------------------------------------------
    //      Регистровые ступени на контролируемом тактовом сигнале
    initial mon_reg = '0;
    always @(posedge reset, posedge monclk)
        if (reset)
            mon_reg <= '0;
        else
            mon_reg <= {mon_reg[CYCLES - 2 : 0], ~ref_reg[CYCLES - 1]};
    
    //------------------------------------------------------------------------------------
    //      Регистровые ступени на опорном тактовом сигнале
    initial ref_reg = '0;
    always @(posedge reset, posedge refclk)
        if (reset)
            ref_reg <= '0;
        else
            ref_reg <= {ref_reg[CYCLES - 2 : 0], mon_reg[CYCLES - 1]};
    
    //------------------------------------------------------------------------------------
    //      Регистр импульсов наличия контролируемого тактового сигнала
    initial pulse_reg ='0;
    always @(posedge reset, posedge refclk)
        if (reset)
            pulse_reg <= '0;
        else
            pulse_reg <= ref_reg[CYCLES - 2] ^ ref_reg[CYCLES - 1];
    
    //------------------------------------------------------------------------------------
    //      Счетчик обнаружения
    initial detect_cnt = CMAX;
    always @(posedge reset, posedge refclk)
        if (reset)
            detect_cnt <= CMAX;
        else if (pulse_reg)
            detect_cnt <= '0;
        else if (detect_cnt == CMAX)
            detect_cnt <= detect_cnt;
        else
            detect_cnt <= detect_cnt + 1'b1;
    
    //------------------------------------------------------------------------------------
    //      Регистр обнаружения
    initial detect_reg = '0;
    always @(posedge reset, posedge refclk)
        if (reset)
            detect_reg <= '0;
        else
            detect_reg <= ~(detect_cnt == CMAX);
    assign detected = detect_reg;
    
endmodule: clockmon