module iterated_fixed_to_float_tb ();
    
    //------------------------------------------------------------------------------------
    //      Описание констант
    localparam              WIDTH = 8;  // Разрядность входных данных (знакового целого)
    
    //------------------------------------------------------------------------------------
    //      Описание сигналов
    logic                   reset;
    logic                   clk;
    //
    logic                   start;
    logic                   ready;
    logic                   done;
    //
    logic [WIDTH - 1 : 0]   fixed;
    logic [31 : 0]          float;
    shortreal               res;
    
    //------------------------------------------------------------------------------------
    //      Сброс
    initial begin
        #00 reset = '1;
        #15 reset = '0;
    end
    
    //------------------------------------------------------------------------------------
    //      Тактирование
    initial clk = '1;
    always  clk = #05 ~clk;
    
    //------------------------------------------------------------------------------------
    //      Инициализация
    initial begin
        start = 0;
        fixed = 0;
    end
    
    //------------------------------------------------------------------------------------
    //      Модуль итерационного перевода знакового целого произвольной разрядности
    //      в число с плавающей точкой одинарной точности
    iterated_fixed_to_float
    #(
        .WIDTH      (WIDTH)     // Разрядность входных данных (знакового целого)
    )
    the_iterated_fixed_to_float
    (
        // Сброс и тактирование
        .reset      (reset),    // i
        .clk        (clk),      // i
        
        // Интерфейс управления
        .start      (start),    // i
        .ready      (ready),    // o
        .done       (done),     // o
        
        // Интерфейс входных данных
        .fixed      (fixed),    // i  [WIDTH - 1 : 0]
        
        // Интерфейс выходных данных
        .float      (float)     // o  [31 : 0]
    ); // the_iterated_fixed_to_float
    
    //------------------------------------------------------------------------------------
    //      Результат в формате с плавающей точкой
    assign res = $bitstoshortreal(float);
    
    //------------------------------------------------------------------------------------
    //      Тестирование
    initial begin
        #100;
        @(posedge clk);
        start = 1;
        while(1) begin
            @(posedge clk);
            while(~ready) @(posedge clk);
            fixed++;
        end
    end
    
endmodule // iterated_fixed_to_float_tb