/*
    //------------------------------------------------------------------------------------
    //      ������������� ���������� ���������� DataStream
    //      (��������� ��������������)
    ds_mux
    #(
        .WIDTH      (), // ����������� ������
        .INPUTS     ()  // ���������� ������� ����������� (����� 1-��)
    )
    the_ds_mux
    (
        // ����� � ������������
        .reset      (), // i  �� ������������
        .clk        (), // i  �� ������������
        
        // ���� ������ ��������� �����
        .select     (), // i  [$clog2(INPUTS) - 1 : 0]
        
        // ������� ��������� ����������
        .i_dat      (), // i  [INPUTS - 1 : 0][WIDTH - 1 : 0]
        .i_val      (), // i  [INPUTS - 1 : 0]
        .i_rdy      (), // o  [INPUTS - 1 : 0]
        
        // �������� ��������� ���������
        .o_dat      (), // o  [WIDTH - 1 : 0]
        .o_val      (), // o
        .o_rdy      ()  // i
    ); // the_ds_mux
*/

module ds_mux
#(
    parameter int unsigned                          WIDTH   = 8,    // ����������� ������
    parameter int unsigned                          INPUTS  = 2     // ���������� ������� ����������� (����� 1-��)
)
(
    // ����� � ������������
    input  logic                                    reset,          // �� ������������
    input  logic                                    clk,            // �� ������������
    
    // ���� ������ ��������� �����
    input  logic [$clog2(INPUTS) - 1 : 0]           select,
    
    // ������� ��������� ����������
    input  logic [INPUTS - 1 : 0][WIDTH - 1 : 0]    i_dat,
    input  logic [INPUTS - 1 : 0]                   i_val,
    output logic [INPUTS - 1 : 0]                   i_rdy,
    
    // �������� ��������� ���������
    output logic [WIDTH - 1 : 0]                    o_dat,
    output logic                                    o_val,
    input  logic                                    o_rdy
);
    //------------------------------------------------------------------------------------
    //      �������� ��������
    logic [INPUTS - 1 : 0]                          select_pos;
    
    //------------------------------------------------------------------------------------
    //      ����������� ��� ����������� ������
    always_comb begin
        select_pos = {INPUTS{1'b0}};
        select_pos[select] = 1'b1;
    end
    
    //------------------------------------------------------------------------------------
    //      ������������ �������� ���������� ��������� ������� �����������
    assign i_rdy = select_pos & {INPUTS{o_rdy}};
    
    //------------------------------------------------------------------------------------
    //      ������������ �������� ��������� ���������� ����������
    assign o_dat = i_dat[select];
    assign o_val = i_val[select];
    
endmodule // ds_mux