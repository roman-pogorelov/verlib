/*
    //------------------------------------------------------------------------------------
    //      Арбитр доступа нескольких абонентов к одному ресурсу
    arbitrator
    #(
        .REQS           (), // Количество абонентов (REQS > 1)
        .SCHEME         ()  // Схема арбитража ("RR" - циклическая, "FP" - фиксированная)
    )
    the_arbitrator
    (
        // Сброс и тактирование
        .reset          (), // i
        .clk            (), // i
        
        // Вектор запросов на обслуживание
        .req            (), // i  [REQS - 1 : 0]
        
        // Готовность обработать запрос
        .rdy            (), // i
        
        // Вектор гранта на обслуживание
        .gnt            (), // o  [REQS - 1 : 0]
        
        // Номер порта, получившего грант
        .num            ()  // o  [$clog2(REQS) - 1 : 0]
    ); // the_arbitrator
*/

module arbitrator
#(
    parameter                           REQS    = 4,    // Количество абонентов (REQS > 1)
    parameter                           SCHEME  = "FP"  // Схема арбитража ("RR" - циклическая, "FP" - фиксированная)
)
(
    // Сброс и тактирование
    input  logic                        reset,
    input  logic                        clk,
    
    // Вектор запросов на обслуживание
    input  logic [REQS - 1 : 0]         req,
    
    // Готовность обработать запрос
    input  logic                        rdy,
    
    // Вектор гранта на обслуживание
    output logic [REQS - 1 : 0]         gnt,
    
    // Номер порта, получившего грант
    output logic [$clog2(REQS) - 1 : 0] num
);
    //------------------------------------------------------------------------------------
    //      Описание сигналов
    logic [REQS - 1 : 0]                top_priority;       // Позиция наивысшего приоритета
    logic [REQS - 1 : 0]                top_priority_reg;   // Регистр позиции наивысшего приоритета
    logic [2*REQS - 1 : 0]              gnt_double;         // Вектор "сдвоенного" гранта
    logic [REQS - 1 : 0]                act_gnt;            // "Активный" грант (формируемый исходя из вектора запросов и схемы арбитража)
    logic [REQS - 1 : 0]                pnd_gnt_reg;        // Регистр гранта, ожидающего обслуживания
    logic                               pnd_req_reg;        // Регистр признака необработанного запроса
    
    //------------------------------------------------------------------------------------
    //      Выбор схемы арбитража
    generate
        // Циклическая схема (round-robin)
        if (SCHEME == "RR")
            assign top_priority = top_priority_reg;
        // Фиксированная схема (fixed priority)
        else
            assign top_priority = {{(REQS - 1){1'b0}}, 1'b1};
    endgenerate
    
    //------------------------------------------------------------------------------------
    //      Регистр позиции наивысшего приоритета
    always @(posedge reset, posedge clk)
        if (reset)
            top_priority_reg <= {{(REQS - 1){1'b0}}, 1'b1};
        else if (|req & rdy)
            top_priority_reg <= {gnt[REQS - 2 : 0], gnt[REQS - 1]};
        else
            top_priority_reg <= top_priority_reg;
    
    //------------------------------------------------------------------------------------
    //      Вектор "сдвоенного" гранта
    assign gnt_double = {req, req} & ({~req, ~req} + {{REQS{1'b0}}, top_priority});
    
    //------------------------------------------------------------------------------------
    //      "Активный" грант (формируемый исходя из вектора запросов и схемы арбитража)
    assign act_gnt = gnt_double[2*REQS - 1 : REQS] | gnt_double[REQS - 1 : 0];
    
    //------------------------------------------------------------------------------------
    //      Регистр гранта, ожидающего обслуживания
    always @(posedge reset, posedge clk)
        if (reset)
            pnd_gnt_reg <= '0;
        else if (~pnd_req_reg & |req & ~rdy)
            pnd_gnt_reg <= act_gnt;
        else
            pnd_gnt_reg <= pnd_gnt_reg;
    
    //------------------------------------------------------------------------------------
    //      Регистр признака необработанного запроса
    always @(posedge reset, posedge clk)
        if (reset)
            pnd_req_reg <= '0;
        else if (pnd_req_reg)
            pnd_req_reg <= ~rdy;
        else
            pnd_req_reg <= |req & ~rdy;
    
    //------------------------------------------------------------------------------------
    //      Вектор гранта на обслуживание
    assign gnt = pnd_req_reg ? pnd_gnt_reg : act_gnt;
    
    //------------------------------------------------------------------------------------
    //      Преобразователь позиционного кода в двоичный
    onehot2binary
    #(
        .WIDTH      (REQS)  // Разрядность входа позиционного кода
    )
    gnt2num_conv
    (
        .onehot     (gnt),  // i  [WIDTH - 1 : 0]
        .binary     (num)   // o  [$clog2(WIDTH) - 1 : 0]
    ); // gnt2num_conv
    
endmodule // arbitrator