`ifndef _CORDIC_DEFINES_H_
`define _CORDIC_DEFINES_H_

    // Коэффициент усиления
    localparam logic [63 : 0] CORDIC_GAIN = 64'h4DBA76D421AF2D34;

    // Таблица элементарных углов поворота
    localparam logic [63 : 0][63 : 0] CORDIC_LUT =
    {
            64'h0000000000000001,
            64'h0000000000000001,
            64'h0000000000000003,
            64'h0000000000000005,
            64'h000000000000000A,
            64'h0000000000000014,
            64'h0000000000000029,
            64'h0000000000000051,
            64'h00000000000000A3,
            64'h0000000000000146,
            64'h000000000000028C,
            64'h0000000000000518,
            64'h0000000000000A30,
            64'h000000000000145F,
            64'h00000000000028BE,
            64'h000000000000517D,
            64'h000000000000A2FA,
            64'h00000000000145F3,
            64'h0000000000028BE6,
            64'h00000000000517CC,
            64'h00000000000A2F98,
            64'h0000000000145F30,
            64'h000000000028BE61,
            64'h0000000000517CC2,
            64'h0000000000A2F983,
            64'h000000000145F307,
            64'h00000000028BE60E,
            64'h000000000517CC1B,
            64'h000000000A2F9837,
            64'h00000000145F306E,
            64'h0000000028BE60DC,
            64'h00000000517CC1B7,
            64'h00000000A2F9836E,
            64'h0000000145F306DD,
            64'h000000028BE60DB9,
            64'h0000000517CC1B72,
            64'h0000000A2F9836E5,
            64'h000000145F306DCA,
            64'h00000028BE60DB94,
            64'h000000517CC1B727,
            64'h000000A2F9836E4E,
            64'h00000145F306DC9D,
            64'h0000028BE60DB939,
            64'h00000517CC1B7270,
            64'h00000A2F9836E4D7,
            64'h0000145F306DC95C,
            64'h000028BE60DB902C,
            64'h0000517CC1B70BF8,
            64'h0000A2F9836D74F7,
            64'h000145F306D5D223,
            64'h00028BE60D82E5E5,
            64'h000517CC19BFD8C3,
            64'h000A2F982950196E,
            64'h00145F30012374F7,
            64'h0028BE5D7661566F,
            64'h00517CA68DA1866E,
            64'h00A2F8AA23A8855D,
            64'h0145EC3CB8504C53,
            64'h028BAFC2B208C4F1,
            64'h05161A861CB135DA,
            64'h0A2223A83BBB3437,
            64'h13F670B6BDC73D1C,
            64'h25C80A3B3BE610CD,
            64'h4000000000000000
    };

`endif // _CORDIC_DEFINES_H_