`timescale  1ns / 1ps
module alt_rom_sin_cos_tb ();
    
    //------------------------------------------------------------------------------------
    //      Описание констант
    localparam int unsigned WIDTH   = 16;               // Разрядность
    parameter               HEXFILE = "sin-lut.hex";    // HEX-файл с предварительно расчитанный таблицей синусов

    //------------------------------------------------------------------------------------
    //      Объявление сигналов
    logic                   reset;
    logic                   clk;
    logic                   clkena;
    logic [WIDTH - 1 : 0]   arg;
    logic [WIDTH - 1 : 0]   sin;
    logic [WIDTH - 1 : 0]   cos;
    
    //------------------------------------------------------------------------------------
    //      Сброс
    initial begin
        #00 reset = '1;
        #15 reset = '0;
    end
    
    //------------------------------------------------------------------------------------
    //      Тактирование
    initial clk = '1;
    always  clk = #05 ~clk;
    
    //------------------------------------------------------------------------------------
    //      Инициализация
    initial begin
        clkena  = 1;
        arg     = 0;
    end
    
    //------------------------------------------------------------------------------------
    //      Модуль табличного вычисления значений функций sin(x) и cos(x)
    alt_rom_sin_cos
    #(
        .WIDTH      (WIDTH),    // Разрядность
        .HEXFILE    (HEXFILE)   // HEX-файл с предварительно расчитанный таблицей синусов
    )
    the_alt_rom_sin_cos
    (
        // Сброс и тактирование
        .reset      (reset),    // i
        .clk        (clk),      // i
        
        // Разрешение тактирования
        .clkena     (clkena),   // i
        
        // Значение аргумента
        .arg        (arg),      // i  [WIDTH - 1 : 0]
        
        // Значения sin(arg), cos(arg)
        .sin        (sin),      // o  [WIDTH - 1 : 0]
        .cos        (cos)       // o  [WIDTH - 1 : 0]
    ); // the_alt_rom_sin_cos
    
    //------------------------------------------------------------------------------------
    //      Тестирование
    initial begin
        #100;
        while(1) begin
            @(posedge clk);
            arg = arg + clkena;
        end
    end
    
endmodule: alt_rom_sin_cos_tb
